`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.10.2025 21:36:00
// Design Name: 
// Module Name: time_core
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//// File: time_core.v
module time_core(
        input clk,
        input rst,
        input load_settings,       
        input [5:0] load_sec,
        input [5:0] load_min,
        input [4:0] load_hour,
        input [4:0] load_day,
        input [3:0] load_month,
        output [3:0] actual_month,
        output [4:0] actual_day, actual_hour,
        output [5:0] actual_min, actual_sec,       
        output [7:0] segm,   
        output [7:0] dign,
        output [5:0] led
    );
    
    wire [5:0] sec, min, l;
    wire [4:0] hour; // 5 bit az �r�nak (0-23)
    wire [3:0] month; // 4 bit a h�napnak (1-12)
    wire [31:0] hex;
    wire [7:0] seg, dig;
    wire day_ce, hour_ce, min_ce, sec_ce;
    wire [3:0] mot, mou, dt, du, ht, hu, mit, miu;
      
    // 1Hz enged�ly jel
    wire ce;
    rategen rategenerator(.clk(clk), .rst(rst), .cy(ce));
    
    // m�sodperc sz�ml�l� 0-59, alaphelyzet 0
    bcd_unit_counter #(0, 59, 0) counter_sec (
        .clk(clk), 
        .rst(rst), 
        .ce(ce),
        .load_en(load_settings),
        .load_data(load_sec),
        .q(sec), 
        .cout(sec_ce)
    );
    
    
    // perc sz�ml�l� 0-59, alaphelyzet 20
    bcd_unit_counter #(0, 59, 20) counter_min (
        .clk(clk), 
        .rst(rst), 
        .ce(ce&sec_ce),
        .load_en(load_settings),
        .load_data(load_min),
        .q(min), 
        .cout(min_ce)
    );        
        
        
    // �ra sz�ml�l� 0-23, alaphelyzet 4
   bcd_unit_counter #(0, 23, 4) counter_hour (
        .clk(clk), 
        .rst(rst), 
        .ce(ce&sec_ce&min_ce),
        .load_en(load_settings),
        .load_data({1'b0, load_hour}), // 5 bit a 6 bites portra
        .q(hour), 
        .cout(hour_ce)
    );
  
    
    // nap sz�ml�l� 1-31 h�napt�l f�gg, alaphelyzet 17
    day_counter day_counter (
        .clk(clk),
        .rst(rst),
        .ce(ce&sec_ce&min_ce&hour_ce),
        .load_en(load_settings),
        .load_day(load_day),
        .month_tens(mot),
        .month_units(mou),
        .du(du),
        .dt(dt),
        .cout(day_ce)
    );
    
    
    // h�nap sz�ml�l� 1-12, alaphelyzet 8
     bcd_unit_counter #(1, 12, 8) counter_month (
        .clk(clk), 
        .rst(rst), 
        .ce(ce&sec_ce&min_ce&hour_ce&day_ce),
        .load_en(load_settings),
        .load_data({2'b0, load_month}), // 4 bit a 6 bites portra
        .q(month), 
        .cout()
    );
    
    
    // kijelz� meghajt�
    hex7seg segdecoder ( 
        .val(hex), 
        .cclk(clk), 
        .rst(rst), 
        .seg(seg), 
        .dig(dig)
    );
    
    // led kapcsol�s
    hexled seconds_display (
        .val(sec),
        .rst(rst),
        .led(l)    
    );
    
    // segmensek l�trehoz�sa sz�mokb�l, t�zesekre �s egyesekre bont�s
    assign miu = min % 10;
    assign mit = min / 10;
    assign hu = hour % 10;
    assign ht = hour / 10;
    assign mou = month % 10;
    assign mot = month / 10;
    
    assign actual_month = month;
    assign actual_day   = dt * 10 + du;
    assign actual_hour  = hour;
    assign actual_min   = min;
    assign actual_sec  = sec;
    
    assign hex = { mot, mou, dt, du, ht, hu, mit, miu };
    assign segm = seg;
    assign dign = ~dig; 
    assign led = l;

endmodule